`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module c6288_tb ;

reg N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,
      N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,
      N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,
      N511,N528;

reg [2:0]score;

wire N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,
       N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,
       N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,
       N6287,N6288;
	   
c6288 uut(.gat1(N1),.gat18(N18),.gat35(N35),.gat52(N52),.gat69(N69),.gat86(N86),.gat103(N103),.gat120(N120),.gat137(N137),.gat154(N154),.gat171(N171),.gat188(N188),.gat205(N205),.gat222(N222),.gat239(N239),.gat256(N256),.gat273(N273),.gat290(N290),.gat307(N307),.gat324(N324),.gat341(N341),.gat358(N358),.gat375(N375),.gat392(N392),.gat409(N409),.gat426(N426),.gat443(N443),.gat460(N460),.gat477(N477),.gat494(N494),.gat511(N511),.gat528(N528),.gat_out545(N545),.gat_out1581(N1581),.gat_out1901(N1901),.gat_out2223(N2223),.gat_out2548(N2548),.gat_out2877(N2877),.gat_out3211(N3211),.gat_out3552(N3552),.gat_out3895(N3895),.gat_out4241(N4241),.gat_out4591(N4591),.gat_out4946(N4946),.gat_out5308(N5308),.gat_out5672(N5672),.gat_out5971(N5971),.gat_out6123(N6123),.gat_out6150(N6150),.gat_out6160(N6160),.gat_out6170(N6170),.gat_out6180(N6180),.gat_out6190(N6190),.gat_out6200(N6200),.gat_out6210(N6210),.gat_out6220(N6220),.gat_out6230(N6230),.gat_out6240(N6240),.gat_out6250(N6250),.gat_out6260(N6260),.gat_out6270(N6270),.gat_out6280(N6280),.gat_out6287(N6287),.gat_out6288(N6288));

initial begin


score <= 3'b000;

//111110000011111000001111100000111110//
N1 <= 1; N18 <= 1 ; N35 <= 1 ; N52 <= 0 ; N69 <= 0 ; N86 <= 0 ; N103 <= 0 ; N120 <= 0 ; N137 <= 0 ; N154 <= 0 ; N171 <= 0 ; N188 <= 0 ; N205 <= 1 ; N222 <= 1 ; N239 <= 1 ; N256 <= 1 ; N273 <= 1 ; N290 <= 0 ; N307 <= 0 ; N324 <= 0 ; N341 <= 0 ; N358 <= 1 ; N375 <= 1 ; N392 <= 1 ; N409 <= 1 ; N426 <= 1 ; N443 <= 1 ; N460 <= 1 ; N477 <= 1 ; N494 <= 0 ; N511 <= 0 ; N528 <= 0 ; 
#10
$display(" input pattern = ",N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528 ," --> golden value = 11100100111100111100011110111000 "); 
$display(" your answer = " ,N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288); 
if (N545 == 1'b1 && N1581 == 1'b1 && N1901 == 1'b1 && N2223 == 1'b0 && N2548 == 1'b0 && N2877 == 1'b1 && N3211 == 1'b0 && N3552 == 1'b0 && N3895 == 1'b1 && N4241 == 1'b1 && N4591 == 1'b1 && N4946 == 1'b1 && N5308 == 1'b0 && N5672 == 1'b0 && N5971 == 1'b1 && N6123 == 1'b1 && N6150 == 1'b1 && N6160 == 1'b1 && N6170 == 1'b0 && N6180 == 1'b0 && N6190 == 1'b0 && N6200 == 1'b1 && N6210 == 1'b1 && N6220 == 1'b1 && N6230 == 1'b1 && N6240 == 1'b0 && N6250 == 1'b1 && N6260 == 1'b1 && N6270 == 1'b1 && N6280 == 1'b0 && N6287 == 1'b0 && N6288 == 1'b0)
begin
	score = score + 3'b001;
end
//110011111111111111110000000000001100//
N1 <= 1; N18 <= 1 ; N35 <= 1 ; N52 <= 1 ; N69 <= 1 ; N86 <= 1 ; N103 <= 1 ; N120 <= 1 ; N137 <= 1 ; N154 <= 1 ; N171 <= 1 ; N188 <= 1 ; N205 <= 1 ; N222 <= 1 ; N239 <= 1 ; N256 <= 1 ; N273 <= 1 ; N290 <= 1 ; N307 <= 1 ; N324 <= 1 ; N341 <= 1 ; N358 <= 1 ; N375 <= 1 ; N392 <= 1 ; N409 <= 1 ; N426 <= 1 ; N443 <= 1 ; N460 <= 1 ; N477 <= 1 ; N494 <= 1 ; N511 <= 1 ; N528 <= 1 ; 
#10
$display(" input pattern = ",N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528 ," --> golden value = 10000000000000000111111111111111 "); 
$display(" your answer = " , N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288); 
if (N545 == 1'b1 && N1581 == 1'b0 && N1901 == 1'b0 && N2223 == 1'b0 && N2548 == 1'b0 && N2877 == 1'b0 && N3211 == 1'b0 && N3552 == 1'b0 && N3895 == 1'b0 && N4241 == 1'b0 && N4591 == 1'b0 && N4946 == 1'b0 && N5308 == 1'b0 && N5672 == 1'b0 && N5971 == 1'b0 && N6123 == 1'b0 && N6150 == 1'b0 && N6160 == 1'b1 && N6170 == 1'b1 && N6180 == 1'b1 && N6190 == 1'b1 && N6200 == 1'b1 && N6210 == 1'b1 && N6220 == 1'b1 && N6230 == 1'b1 && N6240 == 1'b1 && N6250 == 1'b1 && N6260 == 1'b1 && N6270 == 1'b1 && N6280 == 1'b1 && N6287 == 1'b1 && N6288 == 1'b1)
begin
	score = score + 3'b001;
end
//000001111111111111110000000000000000//
N1 <= 0; N18 <= 0 ; N35 <= 0 ; N52 <= 0 ; N69 <= 0 ; N86 <= 0 ; N103 <= 0 ; N120 <= 0 ; N137 <= 0 ; N154 <= 0 ; N171 <= 0 ; N188 <= 0 ; N205 <= 0 ; N222 <= 0 ; N239 <= 0 ; N256 <= 0 ; N273 <= 0 ; N290 <= 0 ; N307 <= 0 ; N324 <= 0 ; N341 <= 0 ; N358 <= 0 ; N375 <= 0 ; N392 <= 0 ; N409 <= 0 ; N426 <= 0 ; N443 <= 0 ; N460 <= 0 ; N477 <= 0 ; N494 <= 0 ; N511 <= 0 ; N528 <= 0 ; 
#10
$display(" input pattern = ",N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528 ," --> golden value = 00000000000000000000000000000000 "); 
$display(" your answer = " , N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288); 
if (N545 == 1'b0 && N1581 == 1'b0 && N1901 == 1'b0 && N2223 == 1'b0 && N2548 == 1'b0 && N2877 == 1'b0 && N3211 == 1'b0 && N3552 == 1'b0 && N3895 == 1'b0 && N4241 == 1'b0 && N4591 == 1'b0 && N4946 == 1'b0 && N5308 == 1'b0 && N5672 == 1'b0 && N5971 == 1'b0 && N6123 == 1'b0 && N6150 == 1'b0 && N6160 == 1'b0 && N6170 == 1'b0 && N6180 == 1'b0 && N6190 == 1'b0 && N6200 == 1'b0 && N6210 == 1'b0 && N6220 == 1'b0 && N6230 == 1'b0 && N6240 == 1'b0 && N6250 == 1'b0 && N6260 == 1'b0 && N6270 == 1'b0 && N6280 == 1'b0 && N6287 == 1'b0 && N6288 == 1'b0)
begin
	score = score + 3'b001;
end
//000001111111111111110000000000011111//
N1 <= 1; N18 <= 1 ; N35 <= 1 ; N52 <= 0 ; N69 <= 0 ; N86 <= 0 ; N103 <= 0 ; N120 <= 0 ; N137 <= 0 ; N154 <= 0 ; N171 <= 0 ; N188 <= 0 ; N205 <= 0 ; N222 <= 0 ; N239 <= 0 ; N256 <= 0 ; N273 <= 0 ; N290 <= 1 ; N307 <= 1 ; N324 <= 1 ; N341 <= 1 ; N358 <= 0 ; N375 <= 0 ; N392 <= 0 ; N409 <= 0 ; N426 <= 0 ; N443 <= 1 ; N460 <= 1 ; N477 <= 1 ; N494 <= 1 ; N511 <= 1 ; N528 <= 1 ; 
#10
$display(" input pattern = ",N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528 ," --> golden value = 01001011001001110110000000000000 "); 
$display(" your answer = " , N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288); 
if (N545 == 1'b0 && N1581 == 1'b1 && N1901 == 1'b0 && N2223 == 1'b0 && N2548 == 1'b1 && N2877 == 1'b0 && N3211 == 1'b1 && N3552 == 1'b1 && N3895 == 1'b0 && N4241 == 1'b0 && N4591 == 1'b1 && N4946 == 1'b0 && N5308 == 1'b0 && N5672 == 1'b1 && N5971 == 1'b1 && N6123 == 1'b1 && N6150 == 1'b0 && N6160 == 1'b1 && N6170 == 1'b1 && N6180 == 1'b0 && N6190 == 1'b0 && N6200 == 1'b0&& N6210 == 1'b0 && N6220 == 1'b0 && N6230 == 1'b0 && N6240 == 1'b0 && N6250 == 1'b0 && N6260 == 1'b0 && N6270 == 1'b0 && N6280 == 1'b0 && N6287 == 1'b0 && N6288 == 1'b0)
begin
	score = score + 3'b001;
end
//111111111111111111001100000000000000//
N1 <= 0; N18 <= 0 ; N35 <= 0 ; N52 <= 0 ; N69 <= 0 ; N86 <= 1 ; N103 <= 1 ; N120 <= 1 ; N137 <= 1 ; N154 <= 1 ; N171 <= 1 ; N188 <= 1 ; N205 <= 0 ; N222 <= 0 ; N239 <= 0 ; N256 <= 0 ; N273 <= 0 ; N290 <= 0 ; N307 <= 1 ; N324 <= 1 ; N341 <= 1 ; N358 <= 1 ; N375 <= 1 ; N392 <= 1 ; N409 <= 0 ; N426 <= 0 ; N443 <= 0 ; N460 <= 0 ; N477 <= 0 ; N494 <= 0 ; N511 <= 1 ; N528 <= 1 ; 
#10
$display(" input pattern = ",N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528 ," --> golden value = 00000001000001011110111111010000 "); 
$display(" your answer = " , N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288); 
if (N545 == 1'b0 && N1581 == 1'b0 && N1901 == 1'b0 && N2223 == 1'b0 && N2548 == 1'b0 && N2877 == 1'b0 && N3211 == 1'b0 && N3552 == 1'b1 && N3895 == 1'b0 && N4241 == 1'b0 && N4591 == 1'b0&& N4946 == 1'b0 && N5308 == 1'b0 && N5672 == 1'b1 && N5971 == 1'b0 && N6123 == 1'b1 && N6150 == 1'b1 && N6160 == 1'b1 && N6170 == 1'b1 && N6180 == 1'b0 && N6190 == 1'b1 && N6200 == 1'b1 && N6210 == 1'b1 && N6220 == 1'b1 && N6230 == 1'b1 && N6240 == 1'b1 && N6250 == 1'b0 && N6260 == 1'b1 && N6270 == 1'b0 && N6280 == 1'b0 && N6287 == 1'b0 && N6288 == 1'b0)
begin
	score = score + 3'b001;
end
if (score == 3'b101)
begin
$display("You're all correct!!!");
$display("  ***    *** ");
$display(" *****  *****");
$display("**************");
$display(" ************ ");
$display("  **********  ");
$display("   ********   ");
$display("    ******    ");
$display("     ****     ");
$display("      **      ");
end
else
$display("WRONG");

end
  
endmodule